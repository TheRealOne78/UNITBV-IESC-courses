//---------------------------------------------------------------
// Proiect    : Electronica Digitala
//              Carte de invatatura
// Autor      : Dan NICULA 
// An         : 2025
//---------------------------------------------------------------
// Descriere  : Multiplexor 5x1 cu selecție one-hot, data pe 8b
//---------------------------------------------------------------

module mux5x1_8b_onehot (
input      [5   -1 :0] sel      , // selectie, 5 biti, one-hot
input      [8*5 -1 :0] data_in  , // data de intrare, 5 x 8 biti
output reg [8   -1 :0] data_out   // data de iesire, 8 biti
);

// codul aici

endmodule // mux5x1_8b_onehot

