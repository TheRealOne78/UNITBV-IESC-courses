//---------------------------------------------------------------
// Proiect    : Electronica Digitala
//              Carte de invatatura
// Autor      : Dan NICULA 
// An         : 2025
//---------------------------------------------------------------
// Descriere  : Codificator cu prioritate de 8 biti
//---------------------------------------------------------------

module encoder8b (
input   [8 -1:0] data_in  , // data de intrare
output  [3 -1:0] data_out , // data de iesire
output           valid      // data de iesire valida
);

// codul aici

endmodule // encoder8b

