//---------------------------------------------------------------
// Proiect    : Electronica Digitala
//              Carte de invatatura
// Autor      : Dan NICULA 
// An         : 2025
//---------------------------------------------------------------
// Descriere  : Codificator cu prioritate de 8 biti, 
//              codare iesire one-hot
//---------------------------------------------------------------

module encoder8b_onehot (
input   [8 -1:0] data_in  , // data de intrare
output  [8 -1:0] data_out , // data de iesire, codata one-hot
output           valid      // data de iesire valida
);

// codul aici

endmodule // encoder8b_onehot
