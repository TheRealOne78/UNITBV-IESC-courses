//---------------------------------------------------------------
// Proiect    : Electronica Digitala
//              Carte de invatatura
// Autor      : Dan NICULA 
// An         : 2025
//---------------------------------------------------------------
// Descriere  : Generator numerele lui Fibonacci
//---------------------------------------------------------------

///// 10 ////////////////////////////////////////////////////////
module fib  (
input              clk       , // ceas (front pozitiv)
input              rst_n     , // reset asincron activ 0
input              ce        , // chip enable, activ 1
input      [4 : 0] idx       , // index numar, in domeniul 0..19
output reg [? : 0] fib_out     // numarul lui Fibonacci
                               //   asociat indexului idx
);

// codul aici

endmodule   // fib
